`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/21/2024 01:30:20 PM
// Design Name: 
// Module Name: SEQ_STORAGE
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module SEQ_STORAGE(
    input BTN,
    input [7:0] LEDS,
    input CLK,
    output LD,
    output [7:0] SEQ
    );
    
    
    
endmodule
